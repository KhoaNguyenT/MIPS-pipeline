//================================================
//  University  : UIT - www.uit.edu.vn
//  Course name : System-on-Chip Design
//  Lab name    : lab3
//  File name   : rom.v
//  Author      : Pham Thanh Hung
//  Date        : Oct 21, 2017
//  Version     : 1.0
//-------------------------------------------------
// Modification History
//
//================================================
module rom(
//input
addr,
//output
data
);

input [31:0] addr;
output [31:0] data;

reg [31:0] data;
`define ADD 6'b100000
`define SUB 6'b100010
`define OP_0 6'h0
`define LW 6'b100011
//
//reg [31:0] mem [0:1023];
//assign data = mem[addr];
//op-6bit|rd-5bit|rt-5bit|rs-5bit|shamt-5bit|function-6bit|
//ADD R3,R2,R1;
//SUB R4,R3,R7;
//LW  R8,4(R3);

always @(*) begin
    case(addr)
    32'h00000000: data = 32'b00000000000000000000000000000000; //DO NOTHING
    32'h00000004: data = 32'b00000000000000000000000000000000; //DO NOTHING
    32'h00000008: data = 32'b00111100000010000000000000010000; //lui t0 0x10        //0x3C080010
    32'h0000000c: data = 32'b00111100000010010000000000100000; //lui t1 0x20        //0x3C090020
    32'h00000010: data = 32'b00000000000000000000000000000000; //DO NOTHING
    32'h00000014: data = 32'b00000000000000000000000000000000; //DO NOTHING
    32'h00000018: data = 32'b00000000000000000000000000000000; //DO NOTHING
    32'h0000001c: data = 32'b00000001001010000101000000100000; //add t2 t1 t0       //0x01285020
    32'h00000020: data = 32'b00000001001010000101100000100100; //and t3 t1 t0       //0x01285824
    32'h00000024: data = 32'b00000001001010000110000000100101; //or t4 t1 t0        //0x01286025
    32'h00000028: data = 32'b00000001001010000110100000100010; //sub t5 t1 t0       //0x01286822
    32'h0000002c: data = 32'b00000001000010010111000000101010; //slt t6 t0 t1       //0x0109702A
    32'h00000030: data = 32'b00010001000010010000000000000000; //beq t0 t1 0x0      //0x11090000
    32'h00000034: data = 32'b10101101011011000000000000000001; //sw t4 0x1 ($t3)    //0xAD6C0001
    32'h00000038: data = 32'b00100001001000000000000000100000; //addi r0 t1 0x20    //0x21200020
    32'h0000003c: data = 32'b10001101011011110000000000000001; //lw t7 0x1 ($t3)    //0x8D6F0001
    32'h00000040: data = 32'b00010001100010100000000000000000; //beq t4 t2 0x0      //0x118A0000
//    32'h00000040: data = 32'b00000000000000000000000000000000; //DO NOTHING
//    32'h00000044: data = 32'b00000000000000000000000000000000; //DO NOTHING
//    32'h00000048: data = 32'b00000000000000000000000000000000; //DO NOTHING
//    32'h0000004c: data = 32'b00000000000000000000000000000000; //DO NOTHING
//    32'h00000050: data = 32'b00000000000000000000000000000000; //DO NOTHING
    
    //insert your instructions here
    default: data = 32'hFFFF_FFFF;
    endcase

end

endmodule